class ALU_configuration extends uvm_object;
	`uvm_object_utils(ALU_configuration)

	function new(string name = "");
		super.new(name);
	endfunction: new
endclass: ALU_configuration