`ifndef Guard_MACRO
`define Guard_MACRO

`define no_op 3'b000
`define add_op 3'b001
`define and_op 3'b010
`define xor_op 3'b011
`define mul_op 3'b100

`endif